`define SIZE 8