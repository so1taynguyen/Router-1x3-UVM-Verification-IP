package router_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "tb_defs.sv"
    `include "router_trans.sv"
    `include "router_env_config.sv"
    `include "router_drv.sv"
    `include "router_mon.sv"
    `include "router_sequencer.sv"
    `include "router_agent.sv"
    `include "router_scoreboard.sv"
    `include "router_env.sv"
    `include "router_seqs.sv"
    `include "router_test_lib.sv"
    
endpackage